// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MMU::*;

import HostInterface::*;

// generated by tool
import GeneralRequest::*;
import GeneralIndication::*;

`ifndef BSIM
import Xilinx       :: *;
import XilinxCells ::*;
import DefaultValue    :: *;
`endif
import Clocks :: *;


// defined by user
import Main::*;

import AuroraExtImport::*;
import AuroraCommon::*;

typedef enum {GeneralIndicationPortal, GeneralRequestPortal, 
   HostMemServerIndicationPortal, HostMemServerRequestPortal, HostMMURequestPortal, HostMMUIndicationPortal
   } IfcNames deriving (Eq,Bits);

(* synthesize *)
module mkConnectalTop#(Clock clk250, Reset rst250) (ConnectalTop#(PhysAddrWidth,DataBusWidth,AuroraExtPins,NumberOfMasters));

   Clock curClk <- exposeCurrentClock;
   Reset curRst <- exposeCurrentReset;

   GeneralIndicationProxy generalIndicationProxy <- mkGeneralIndicationProxy(GeneralIndicationPortal);

   MainIfc hwmain <- mkMain(generalIndicationProxy.ifc, clk250, rst250);
   GeneralRequestWrapper generalRequestWrapper <- mkGeneralRequestWrapper(GeneralRequestPortal,hwmain.request);

   Vector#(2,StdPortal) portals;
   portals[0] = generalRequestWrapper.portalIfc;
   portals[1] = generalIndicationProxy.portalIfc; 
   
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;

   interface AuroraExtPins pins;
      interface Aurora_Pins aurora_ext = hwmain.aurora_ext;
      interface Aurora_Clock_Pins aurora_quad119 = hwmain.aurora_quad119;
   endinterface
endmodule

export mkConnectalTop;
export AuroraExtPins;

